library ieee;

use ieee.std_logic_1164.all;

entity
  BrentKung
is
port
  ( 
 
    
    a_0 : in std_logic
  ; a_1 : in std_logic
  ; a_2 : in std_logic
  ; a_3 : in std_logic
  ; a_4 : in std_logic
  ; a_5 : in std_logic
  ; a_6 : in std_logic
  ; a_7 : in std_logic
  ; a_8 : in std_logic
  ; a_9 : in std_logic
  ; a_10 : in std_logic
  ; a_11 : in std_logic
  ; a_12 : in std_logic
  ; a_13 : in std_logic
  ; a_14 : in std_logic
  ; a_15 : in std_logic
  ; a_16 : in std_logic
  ; a_17 : in std_logic
  ; a_18 : in std_logic
  ; a_19 : in std_logic
  ; a_20 : in std_logic
  ; a_21 : in std_logic
  ; a_22 : in std_logic
  ; a_23 : in std_logic
  ; a_24 : in std_logic
  ; a_25 : in std_logic
  ; a_26 : in std_logic
  ; a_27 : in std_logic
  ; a_28 : in std_logic
  ; a_29 : in std_logic
  ; a_30 : in std_logic
  ; a_31 : in std_logic
  ; a_32 : in std_logic
  ; a_33 : in std_logic
  ; a_34 : in std_logic
  ; a_35 : in std_logic
  ; a_36 : in std_logic
  ; a_37 : in std_logic
  ; a_38 : in std_logic
  ; a_39 : in std_logic
  ; a_40 : in std_logic
  ; a_41 : in std_logic
  ; a_42 : in std_logic
  ; a_43 : in std_logic
  ; a_44 : in std_logic
  ; a_45 : in std_logic
  ; a_46 : in std_logic
  ; a_47 : in std_logic
  ; a_48 : in std_logic
  ; a_49 : in std_logic
  ; a_50 : in std_logic
  ; a_51 : in std_logic
  ; a_52 : in std_logic
  ; a_53 : in std_logic
  ; a_54 : in std_logic
  ; a_55 : in std_logic
  ; a_56 : in std_logic
  ; a_57 : in std_logic
  ; a_58 : in std_logic
  ; a_59 : in std_logic
  ; a_60 : in std_logic
  ; a_61 : in std_logic
  ; a_62 : in std_logic
  ; a_63 : in std_logic
  ; b_0 : in std_logic
  ; b_1 : in std_logic
  ; b_2 : in std_logic
  ; b_3 : in std_logic
  ; b_4 : in std_logic
  ; b_5 : in std_logic
  ; b_6 : in std_logic
  ; b_7 : in std_logic
  ; b_8 : in std_logic
  ; b_9 : in std_logic
  ; b_10 : in std_logic
  ; b_11 : in std_logic
  ; b_12 : in std_logic
  ; b_13 : in std_logic
  ; b_14 : in std_logic
  ; b_15 : in std_logic
  ; b_16 : in std_logic
  ; b_17 : in std_logic
  ; b_18 : in std_logic
  ; b_19 : in std_logic
  ; b_20 : in std_logic
  ; b_21 : in std_logic
  ; b_22 : in std_logic
  ; b_23 : in std_logic
  ; b_24 : in std_logic
  ; b_25 : in std_logic
  ; b_26 : in std_logic
  ; b_27 : in std_logic
  ; b_28 : in std_logic
  ; b_29 : in std_logic
  ; b_30 : in std_logic
  ; b_31 : in std_logic
  ; b_32 : in std_logic
  ; b_33 : in std_logic
  ; b_34 : in std_logic
  ; b_35 : in std_logic
  ; b_36 : in std_logic
  ; b_37 : in std_logic
  ; b_38 : in std_logic
  ; b_39 : in std_logic
  ; b_40 : in std_logic
  ; b_41 : in std_logic
  ; b_42 : in std_logic
  ; b_43 : in std_logic
  ; b_44 : in std_logic
  ; b_45 : in std_logic
  ; b_46 : in std_logic
  ; b_47 : in std_logic
  ; b_48 : in std_logic
  ; b_49 : in std_logic
  ; b_50 : in std_logic
  ; b_51 : in std_logic
  ; b_52 : in std_logic
  ; b_53 : in std_logic
  ; b_54 : in std_logic
  ; b_55 : in std_logic
  ; b_56 : in std_logic
  ; b_57 : in std_logic
  ; b_58 : in std_logic
  ; b_59 : in std_logic
  ; b_60 : in std_logic
  ; b_61 : in std_logic
  ; b_62 : in std_logic
  ; b_63 : in std_logic

  
  ; sum_0 : out std_logic
  ; sum_1 : out std_logic
  ; sum_2 : out std_logic
  ; sum_3 : out std_logic
  ; sum_4 : out std_logic
  ; sum_5 : out std_logic
  ; sum_6 : out std_logic
  ; sum_7 : out std_logic
  ; sum_8 : out std_logic
  ; sum_9 : out std_logic
  ; sum_10 : out std_logic
  ; sum_11 : out std_logic
  ; sum_12 : out std_logic
  ; sum_13 : out std_logic
  ; sum_14 : out std_logic
  ; sum_15 : out std_logic
  ; sum_16 : out std_logic
  ; sum_17 : out std_logic
  ; sum_18 : out std_logic
  ; sum_19 : out std_logic
  ; sum_20 : out std_logic
  ; sum_21 : out std_logic
  ; sum_22 : out std_logic
  ; sum_23 : out std_logic
  ; sum_24 : out std_logic
  ; sum_25 : out std_logic
  ; sum_26 : out std_logic
  ; sum_27 : out std_logic
  ; sum_28 : out std_logic
  ; sum_29 : out std_logic
  ; sum_30 : out std_logic
  ; sum_31 : out std_logic
  ; sum_32 : out std_logic
  ; sum_33 : out std_logic
  ; sum_34 : out std_logic
  ; sum_35 : out std_logic
  ; sum_36 : out std_logic
  ; sum_37 : out std_logic
  ; sum_38 : out std_logic
  ; sum_39 : out std_logic
  ; sum_40 : out std_logic
  ; sum_41 : out std_logic
  ; sum_42 : out std_logic
  ; sum_43 : out std_logic
  ; sum_44 : out std_logic
  ; sum_45 : out std_logic
  ; sum_46 : out std_logic
  ; sum_47 : out std_logic
  ; sum_48 : out std_logic
  ; sum_49 : out std_logic
  ; sum_50 : out std_logic
  ; sum_51 : out std_logic
  ; sum_52 : out std_logic
  ; sum_53 : out std_logic
  ; sum_54 : out std_logic
  ; sum_55 : out std_logic
  ; sum_56 : out std_logic
  ; sum_57 : out std_logic
  ; sum_58 : out std_logic
  ; sum_59 : out std_logic
  ; sum_60 : out std_logic
  ; sum_61 : out std_logic
  ; sum_62 : out std_logic
  ; sum_63 : out std_logic
  ; cout : out std_logic
  );
end BrentKung;

architecture
  structural
of
  BrentKung
is
  signal w1 : std_logic;
  signal w2 : std_logic;
  signal w3 : std_logic;
  signal w4 : std_logic;
  signal w5 : std_logic;
  signal w6 : std_logic;
  signal w7 : std_logic;
  signal w8 : std_logic;
  signal w9 : std_logic;
  signal w10 : std_logic;
  signal w11 : std_logic;
  signal w12 : std_logic;
  signal w13 : std_logic;
  signal w14 : std_logic;
  signal w15 : std_logic;
  signal w16 : std_logic;
  signal w17 : std_logic;
  signal w18 : std_logic;
  signal w19 : std_logic;
  signal w20 : std_logic;
  signal w21 : std_logic;
  signal w22 : std_logic;
  signal w23 : std_logic;
  signal w24 : std_logic;
  signal w25 : std_logic;
  signal w26 : std_logic;
  signal w27 : std_logic;
  signal w28 : std_logic;
  signal w29 : std_logic;
  signal w30 : std_logic;
  signal w31 : std_logic;
  signal w32 : std_logic;
  signal w33 : std_logic;
  signal w34 : std_logic;
  signal w35 : std_logic;
  signal w36 : std_logic;
  signal w37 : std_logic;
  signal w38 : std_logic;
  signal w39 : std_logic;
  signal w40 : std_logic;
  signal w41 : std_logic;
  signal w42 : std_logic;
  signal w43 : std_logic;
  signal w44 : std_logic;
  signal w45 : std_logic;
  signal w46 : std_logic;
  signal w47 : std_logic;
  signal w48 : std_logic;
  signal w49 : std_logic;
  signal w50 : std_logic;
  signal w51 : std_logic;
  signal w52 : std_logic;
  signal w53 : std_logic;
  signal w54 : std_logic;
  signal w55 : std_logic;
  signal w56 : std_logic;
  signal w57 : std_logic;
  signal w58 : std_logic;
  signal w59 : std_logic;
  signal w60 : std_logic;
  signal w61 : std_logic;
  signal w62 : std_logic;
  signal w63 : std_logic;
  signal w64 : std_logic;
  signal w65 : std_logic;
  signal w66 : std_logic;
  signal w67 : std_logic;
  signal w68 : std_logic;
  signal w69 : std_logic;
  signal w70 : std_logic;
  signal w71 : std_logic;
  signal w72 : std_logic;
  signal w73 : std_logic;
  signal w74 : std_logic;
  signal w75 : std_logic;
  signal w76 : std_logic;
  signal w77 : std_logic;
  signal w78 : std_logic;
  signal w79 : std_logic;
  signal w80 : std_logic;
  signal w81 : std_logic;
  signal w82 : std_logic;
  signal w83 : std_logic;
  signal w84 : std_logic;
  signal w85 : std_logic;
  signal w86 : std_logic;
  signal w87 : std_logic;
  signal w88 : std_logic;
  signal w89 : std_logic;
  signal w90 : std_logic;
  signal w91 : std_logic;
  signal w92 : std_logic;
  signal w93 : std_logic;
  signal w94 : std_logic;
  signal w95 : std_logic;
  signal w96 : std_logic;
  signal w97 : std_logic;
  signal w98 : std_logic;
  signal w99 : std_logic;
  signal w100 : std_logic;
  signal w101 : std_logic;
  signal w102 : std_logic;
  signal w103 : std_logic;
  signal w104 : std_logic;
  signal w105 : std_logic;
  signal w106 : std_logic;
  signal w107 : std_logic;
  signal w108 : std_logic;
  signal w109 : std_logic;
  signal w110 : std_logic;
  signal w111 : std_logic;
  signal w112 : std_logic;
  signal w113 : std_logic;
  signal w114 : std_logic;
  signal w115 : std_logic;
  signal w116 : std_logic;
  signal w117 : std_logic;
  signal w118 : std_logic;
  signal w119 : std_logic;
  signal w120 : std_logic;
  signal w121 : std_logic;
  signal w122 : std_logic;
  signal w123 : std_logic;
  signal w124 : std_logic;
  signal w125 : std_logic;
  signal w126 : std_logic;
  signal w127 : std_logic;
  signal w128 : std_logic;
  signal w129 : std_logic;
  signal w130 : std_logic;
  signal w131 : std_logic;
  signal w132 : std_logic;
  signal w133 : std_logic;
  signal w134 : std_logic;
  signal w135 : std_logic;
  signal w136 : std_logic;
  signal w137 : std_logic;
  signal w138 : std_logic;
  signal w139 : std_logic;
  signal w140 : std_logic;
  signal w141 : std_logic;
  signal w142 : std_logic;
  signal w143 : std_logic;
  signal w144 : std_logic;
  signal w145 : std_logic;
  signal w146 : std_logic;
  signal w147 : std_logic;
  signal w148 : std_logic;
  signal w149 : std_logic;
  signal w150 : std_logic;
  signal w151 : std_logic;
  signal w152 : std_logic;
  signal w153 : std_logic;
  signal w154 : std_logic;
  signal w155 : std_logic;
  signal w156 : std_logic;
  signal w157 : std_logic;
  signal w158 : std_logic;
  signal w159 : std_logic;
  signal w160 : std_logic;
  signal w161 : std_logic;
  signal w162 : std_logic;
  signal w163 : std_logic;
  signal w164 : std_logic;
  signal w165 : std_logic;
  signal w166 : std_logic;
  signal w167 : std_logic;
  signal w168 : std_logic;
  signal w169 : std_logic;
  signal w170 : std_logic;
  signal w171 : std_logic;
  signal w172 : std_logic;
  signal w173 : std_logic;
  signal w174 : std_logic;
  signal w175 : std_logic;
  signal w176 : std_logic;
  signal w177 : std_logic;
  signal w178 : std_logic;
  signal w179 : std_logic;
  signal w180 : std_logic;
  signal w181 : std_logic;
  signal w182 : std_logic;
  signal w183 : std_logic;
  signal w184 : std_logic;
  signal w185 : std_logic;
  signal w186 : std_logic;
  signal w187 : std_logic;
  signal w188 : std_logic;
  signal w189 : std_logic;
  signal w190 : std_logic;
  signal w191 : std_logic;
  signal w192 : std_logic;
  signal w193 : std_logic;
  signal w194 : std_logic;
  signal w195 : std_logic;
  signal w196 : std_logic;
  signal w197 : std_logic;
  signal w198 : std_logic;
  signal w199 : std_logic;
  signal w200 : std_logic;
  signal w201 : std_logic;
  signal w202 : std_logic;
  signal w203 : std_logic;
  signal w204 : std_logic;
  signal w205 : std_logic;
  signal w206 : std_logic;
  signal w207 : std_logic;
  signal w208 : std_logic;
  signal w209 : std_logic;
  signal w210 : std_logic;
  signal w211 : std_logic;
  signal w212 : std_logic;
  signal w213 : std_logic;
  signal w214 : std_logic;
  signal w215 : std_logic;
  signal w216 : std_logic;
  signal w217 : std_logic;
  signal w218 : std_logic;
  signal w219 : std_logic;
  signal w220 : std_logic;
  signal w221 : std_logic;
  signal w222 : std_logic;
  signal w223 : std_logic;
  signal w224 : std_logic;
  signal w225 : std_logic;
  signal w226 : std_logic;
  signal w227 : std_logic;
  signal w228 : std_logic;
  signal w229 : std_logic;
  signal w230 : std_logic;
  signal w231 : std_logic;
  signal w232 : std_logic;
  signal w233 : std_logic;
  signal w234 : std_logic;
  signal w235 : std_logic;
  signal w236 : std_logic;
  signal w237 : std_logic;
  signal w238 : std_logic;
  signal w239 : std_logic;
  signal w240 : std_logic;
  signal w241 : std_logic;
  signal w242 : std_logic;
  signal w243 : std_logic;
  signal w244 : std_logic;
  signal w245 : std_logic;
  signal w246 : std_logic;
  signal w247 : std_logic;
  signal w248 : std_logic;
  signal w249 : std_logic;
  signal w250 : std_logic;
  signal w251 : std_logic;
  signal w252 : std_logic;
  signal w253 : std_logic;
  signal w254 : std_logic;
  signal w255 : std_logic;
  signal w256 : std_logic;
  signal w257 : std_logic;
  signal w258 : std_logic;
  signal w259 : std_logic;
  signal w260 : std_logic;
  signal w261 : std_logic;
  signal w262 : std_logic;
  signal w263 : std_logic;
  signal w264 : std_logic;
  signal w265 : std_logic;
  signal w266 : std_logic;
  signal w267 : std_logic;
  signal w268 : std_logic;
  signal w269 : std_logic;
  signal w270 : std_logic;
  signal w271 : std_logic;
  signal w272 : std_logic;
  signal w273 : std_logic;
  signal w274 : std_logic;
  signal w275 : std_logic;
  signal w276 : std_logic;
  signal w277 : std_logic;
  signal w278 : std_logic;
  signal w279 : std_logic;
  signal w280 : std_logic;
  signal w281 : std_logic;
  signal w282 : std_logic;
  signal w283 : std_logic;
  signal w284 : std_logic;
  signal w285 : std_logic;
  signal w286 : std_logic;
  signal w287 : std_logic;
  signal w288 : std_logic;
  signal w289 : std_logic;
  signal w290 : std_logic;
  signal w291 : std_logic;
  signal w292 : std_logic;
  signal w293 : std_logic;
  signal w294 : std_logic;
  signal w295 : std_logic;
  signal w296 : std_logic;
  signal w297 : std_logic;
  signal w298 : std_logic;
  signal w299 : std_logic;
  signal w300 : std_logic;
  signal w301 : std_logic;
  signal w302 : std_logic;
  signal w303 : std_logic;
  signal w304 : std_logic;
  signal w305 : std_logic;
  signal w306 : std_logic;
  signal w307 : std_logic;
  signal w308 : std_logic;
  signal w309 : std_logic;
  signal w310 : std_logic;
  signal w311 : std_logic;
  signal w312 : std_logic;
  signal w313 : std_logic;
  signal w314 : std_logic;
  signal w315 : std_logic;
  signal w316 : std_logic;
  signal w317 : std_logic;
  signal w318 : std_logic;
  signal w319 : std_logic;
  signal w320 : std_logic;
  signal w321 : std_logic;
  signal w322 : std_logic;
  signal w323 : std_logic;
  signal w324 : std_logic;
  signal w325 : std_logic;
  signal w326 : std_logic;
  signal w327 : std_logic;
  signal w328 : std_logic;
  signal w329 : std_logic;
  signal w330 : std_logic;
  signal w331 : std_logic;
  signal w332 : std_logic;
  signal w333 : std_logic;
  signal w334 : std_logic;
  signal w335 : std_logic;
  signal w336 : std_logic;
  signal w337 : std_logic;
  signal w338 : std_logic;
  signal w339 : std_logic;
  signal w340 : std_logic;
  signal w341 : std_logic;
  signal w342 : std_logic;
  signal w343 : std_logic;
  signal w344 : std_logic;
  signal w345 : std_logic;
  signal w346 : std_logic;
  signal w347 : std_logic;
  signal w348 : std_logic;
  signal w349 : std_logic;
  signal w350 : std_logic;
  signal w351 : std_logic;
  signal w352 : std_logic;
  signal w353 : std_logic;
  signal w354 : std_logic;
  signal w355 : std_logic;
  signal w356 : std_logic;
  signal w357 : std_logic;
  signal w358 : std_logic;
  signal w359 : std_logic;
  signal w360 : std_logic;
  signal w361 : std_logic;
  signal w362 : std_logic;
  signal w363 : std_logic;
  signal w364 : std_logic;
  signal w365 : std_logic;
  signal w366 : std_logic;
  signal w367 : std_logic;
  signal w368 : std_logic;
  signal w369 : std_logic;
  signal w370 : std_logic;
  signal w371 : std_logic;
  signal w372 : std_logic;
  signal w373 : std_logic;
  signal w374 : std_logic;
  signal w375 : std_logic;
  signal w376 : std_logic;
  signal w377 : std_logic;
  signal w378 : std_logic;
  signal w379 : std_logic;
  signal w380 : std_logic;
  signal w381 : std_logic;
  signal w382 : std_logic;
  signal w383 : std_logic;
  signal w384 : std_logic;
  signal w385 : std_logic;
  signal w386 : std_logic;
  signal w387 : std_logic;
  signal w388 : std_logic;
  signal w389 : std_logic;
  signal w390 : std_logic;
  signal w391 : std_logic;
  signal w392 : std_logic;
  signal w393 : std_logic;
  signal w394 : std_logic;
  signal w395 : std_logic;
  signal w396 : std_logic;
  signal w397 : std_logic;
  signal w398 : std_logic;
  signal w399 : std_logic;
  signal w400 : std_logic;
  signal w401 : std_logic;
  signal w402 : std_logic;
  signal w403 : std_logic;
  signal w404 : std_logic;
  signal w405 : std_logic;
  signal w406 : std_logic;
  signal w407 : std_logic;
  signal w408 : std_logic;
  signal w409 : std_logic;
  signal w410 : std_logic;
  signal w411 : std_logic;
  signal w412 : std_logic;
  signal w413 : std_logic;
  signal w414 : std_logic;
  signal w415 : std_logic;
  signal w416 : std_logic;
  signal w417 : std_logic;
  signal w418 : std_logic;
  signal w419 : std_logic;
  signal w420 : std_logic;
  signal w421 : std_logic;
  signal w422 : std_logic;
  signal w423 : std_logic;
  signal w424 : std_logic;
  signal w425 : std_logic;
  signal w426 : std_logic;
  signal w427 : std_logic;
  signal w428 : std_logic;
  signal w429 : std_logic;
  signal w430 : std_logic;
  signal w431 : std_logic;
  signal w432 : std_logic;
  signal w433 : std_logic;
  signal w434 : std_logic;
  signal w435 : std_logic;
  signal w436 : std_logic;
  signal w437 : std_logic;
  signal w438 : std_logic;
  signal w439 : std_logic;
  signal w440 : std_logic;
  signal w441 : std_logic;
  signal w442 : std_logic;
  signal w443 : std_logic;
  signal w444 : std_logic;
  signal w445 : std_logic;
  signal w446 : std_logic;
  signal w447 : std_logic;
  signal w448 : std_logic;
  signal w449 : std_logic;
  signal w450 : std_logic;
  signal w451 : std_logic;
  signal w452 : std_logic;
  signal w453 : std_logic;
  signal w454 : std_logic;
  signal w455 : std_logic;
  signal w456 : std_logic;
  signal w457 : std_logic;
  signal w458 : std_logic;
  signal w459 : std_logic;
  signal w460 : std_logic;
  signal w461 : std_logic;
  signal w462 : std_logic;
  signal w463 : std_logic;
  signal w464 : std_logic;
  signal w465 : std_logic;
  signal w466 : std_logic;
  signal w467 : std_logic;
  signal w468 : std_logic;
  signal w469 : std_logic;
  signal w470 : std_logic;
  signal w471 : std_logic;
  signal w472 : std_logic;
  signal w473 : std_logic;
  signal w474 : std_logic;
  signal w475 : std_logic;
  signal w476 : std_logic;
  signal w477 : std_logic;
  signal w478 : std_logic;
  signal w479 : std_logic;
  signal w480 : std_logic;
  signal w481 : std_logic;
  signal w482 : std_logic;
  signal w483 : std_logic;
  signal w484 : std_logic;
  signal w485 : std_logic;
  signal w486 : std_logic;
  signal w487 : std_logic;
  signal w488 : std_logic;
  signal w489 : std_logic;
  signal w490 : std_logic;
  signal w491 : std_logic;
  signal w492 : std_logic;
  signal w493 : std_logic;
  signal w494 : std_logic;
  signal w495 : std_logic;
  signal w496 : std_logic;
  signal w497 : std_logic;
  signal w498 : std_logic;
  signal w499 : std_logic;
  signal w500 : std_logic;
  signal w501 : std_logic;
  signal w502 : std_logic;
  signal w503 : std_logic;
  signal w504 : std_logic;
  signal w505 : std_logic;
  signal w506 : std_logic;
  signal w507 : std_logic;
  signal w508 : std_logic;
  signal w509 : std_logic;
  signal w510 : std_logic;
  signal w511 : std_logic;
  signal w512 : std_logic;
  signal w513 : std_logic;
  signal w514 : std_logic;
  signal w515 : std_logic;
  signal w516 : std_logic;
  signal w517 : std_logic;
  signal w518 : std_logic;
  signal w519 : std_logic;
  signal w520 : std_logic;
  signal w521 : std_logic;
  signal w522 : std_logic;
  signal w523 : std_logic;
  signal w524 : std_logic;
  signal w525 : std_logic;
  signal w526 : std_logic;
  signal w527 : std_logic;
  signal w528 : std_logic;
  signal w529 : std_logic;
  signal w530 : std_logic;
  signal w531 : std_logic;
  signal w532 : std_logic;
  signal w533 : std_logic;
  signal w534 : std_logic;
  signal w535 : std_logic;
  signal w536 : std_logic;
  signal w537 : std_logic;
  signal w538 : std_logic;
  signal w539 : std_logic;
  signal w540 : std_logic;
  signal w541 : std_logic;
  signal w542 : std_logic;
  signal w543 : std_logic;
  signal w544 : std_logic;
  signal w545 : std_logic;
  signal w546 : std_logic;
  signal w547 : std_logic;
  signal w548 : std_logic;
  signal w549 : std_logic;
  signal w550 : std_logic;
  signal w551 : std_logic;
  signal w552 : std_logic;
  signal w553 : std_logic;
  signal w554 : std_logic;
  signal w555 : std_logic;
  signal w556 : std_logic;
  signal w557 : std_logic;
  signal w558 : std_logic;
  signal w559 : std_logic;
  signal w560 : std_logic;
  signal w561 : std_logic;
  signal w562 : std_logic;
  signal w563 : std_logic;
  signal w564 : std_logic;
  signal w565 : std_logic;
  signal w566 : std_logic;
  signal w567 : std_logic;
  signal w568 : std_logic;
  signal w569 : std_logic;
  signal w570 : std_logic;
  signal w571 : std_logic;
  signal w572 : std_logic;
  signal w573 : std_logic;
  signal w574 : std_logic;
  signal w575 : std_logic;
  signal w576 : std_logic;
  signal w577 : std_logic;
  signal w578 : std_logic;
  signal w579 : std_logic;
  signal w580 : std_logic;
  signal w581 : std_logic;
  signal w582 : std_logic;
  signal w583 : std_logic;
  signal w584 : std_logic;
  signal w585 : std_logic;
  signal w586 : std_logic;
  signal w587 : std_logic;
  signal w588 : std_logic;
  signal w589 : std_logic;
  signal w590 : std_logic;
  signal w591 : std_logic;
  signal w592 : std_logic;
  signal w593 : std_logic;
  signal w594 : std_logic;
  signal w595 : std_logic;
  signal w596 : std_logic;
  signal w597 : std_logic;
  signal w598 : std_logic;
  signal w599 : std_logic;
  signal w600 : std_logic;
  signal w601 : std_logic;
  signal w602 : std_logic;
  signal w603 : std_logic;
  signal w604 : std_logic;
  signal w605 : std_logic;
  signal w606 : std_logic;
  signal w607 : std_logic;
  signal w608 : std_logic;
  signal w609 : std_logic;
  signal w610 : std_logic;
  signal w611 : std_logic;
  signal w612 : std_logic;
  signal w613 : std_logic;
  signal w614 : std_logic;
  signal w615 : std_logic;
  signal w616 : std_logic;
begin
  c_w2      : entity work.wire  port map (a_0, w2);
  c_w3      : entity work.wire  port map (b_0, w3);
  c_w1      : entity work.xorG  port map (w2, w3, w1);
  c_w6      : entity work.wire  port map (a_1, w6);
  c_w7      : entity work.wire  port map (b_1, w7);
  c_w5      : entity work.xorG  port map (w6, w7, w5);
  c_w8      : entity work.andG  port map (w2, w3, w8);
  c_w4      : entity work.xorG  port map (w5, w8, w4);
  c_w11     : entity work.wire  port map (a_2, w11);
  c_w12     : entity work.wire  port map (b_2, w12);
  c_w10     : entity work.xorG  port map (w11, w12, w10);
  c_w14     : entity work.andG  port map (w6, w7, w14);
  c_w15     : entity work.andG  port map (w5, w8, w15);
  c_w13     : entity work.orG   port map (w14, w15, w13);
  c_w9      : entity work.xorG  port map (w10, w13, w9);
  c_w18     : entity work.wire  port map (a_3, w18);
  c_w19     : entity work.wire  port map (b_3, w19);
  c_w17     : entity work.xorG  port map (w18, w19, w17);
  c_w21     : entity work.andG  port map (w11, w12, w21);
  c_w22     : entity work.andG  port map (w10, w13, w22);
  c_w20     : entity work.orG   port map (w21, w22, w20);
  c_w16     : entity work.xorG  port map (w17, w20, w16);
  c_w25     : entity work.wire  port map (a_4, w25);
  c_w26     : entity work.wire  port map (b_4, w26);
  c_w24     : entity work.xorG  port map (w25, w26, w24);
  c_w29     : entity work.andG  port map (w18, w19, w29);
  c_w30     : entity work.andG  port map (w17, w21, w30);
  c_w28     : entity work.orG   port map (w29, w30, w28);
  c_w32     : entity work.andG  port map (w17, w10, w32);
  c_w31     : entity work.andG  port map (w32, w13, w31);
  c_w27     : entity work.orG   port map (w28, w31, w27);
  c_w23     : entity work.xorG  port map (w24, w27, w23);
  c_w35     : entity work.wire  port map (a_5, w35);
  c_w36     : entity work.wire  port map (b_5, w36);
  c_w34     : entity work.xorG  port map (w35, w36, w34);
  c_w38     : entity work.andG  port map (w25, w26, w38);
  c_w39     : entity work.andG  port map (w24, w27, w39);
  c_w37     : entity work.orG   port map (w38, w39, w37);
  c_w33     : entity work.xorG  port map (w34, w37, w33);
  c_w42     : entity work.wire  port map (a_6, w42);
  c_w43     : entity work.wire  port map (b_6, w43);
  c_w41     : entity work.xorG  port map (w42, w43, w41);
  c_w46     : entity work.andG  port map (w35, w36, w46);
  c_w47     : entity work.andG  port map (w34, w38, w47);
  c_w45     : entity work.orG   port map (w46, w47, w45);
  c_w49     : entity work.andG  port map (w34, w24, w49);
  c_w48     : entity work.andG  port map (w49, w27, w48);
  c_w44     : entity work.orG   port map (w45, w48, w44);
  c_w40     : entity work.xorG  port map (w41, w44, w40);
  c_w52     : entity work.wire  port map (a_7, w52);
  c_w53     : entity work.wire  port map (b_7, w53);
  c_w51     : entity work.xorG  port map (w52, w53, w51);
  c_w55     : entity work.andG  port map (w42, w43, w55);
  c_w56     : entity work.andG  port map (w41, w44, w56);
  c_w54     : entity work.orG   port map (w55, w56, w54);
  c_w50     : entity work.xorG  port map (w51, w54, w50);
  c_w59     : entity work.wire  port map (a_8, w59);
  c_w60     : entity work.wire  port map (b_8, w60);
  c_w58     : entity work.xorG  port map (w59, w60, w58);
  c_w64     : entity work.andG  port map (w52, w53, w64);
  c_w65     : entity work.andG  port map (w51, w55, w65);
  c_w63     : entity work.orG   port map (w64, w65, w63);
  c_w67     : entity work.andG  port map (w51, w41, w67);
  c_w66     : entity work.andG  port map (w67, w45, w66);
  c_w62     : entity work.orG   port map (w63, w66, w62);
  c_w69     : entity work.andG  port map (w67, w49, w69);
  c_w68     : entity work.andG  port map (w69, w27, w68);
  c_w61     : entity work.orG   port map (w62, w68, w61);
  c_w57     : entity work.xorG  port map (w58, w61, w57);
  c_w72     : entity work.wire  port map (a_9, w72);
  c_w73     : entity work.wire  port map (b_9, w73);
  c_w71     : entity work.xorG  port map (w72, w73, w71);
  c_w75     : entity work.andG  port map (w59, w60, w75);
  c_w76     : entity work.andG  port map (w58, w61, w76);
  c_w74     : entity work.orG   port map (w75, w76, w74);
  c_w70     : entity work.xorG  port map (w71, w74, w70);
  c_w79     : entity work.wire  port map (a_10, w79);
  c_w80     : entity work.wire  port map (b_10, w80);
  c_w78     : entity work.xorG  port map (w79, w80, w78);
  c_w83     : entity work.andG  port map (w72, w73, w83);
  c_w84     : entity work.andG  port map (w71, w75, w84);
  c_w82     : entity work.orG   port map (w83, w84, w82);
  c_w86     : entity work.andG  port map (w71, w58, w86);
  c_w85     : entity work.andG  port map (w86, w61, w85);
  c_w81     : entity work.orG   port map (w82, w85, w81);
  c_w77     : entity work.xorG  port map (w78, w81, w77);
  c_w89     : entity work.wire  port map (a_11, w89);
  c_w90     : entity work.wire  port map (b_11, w90);
  c_w88     : entity work.xorG  port map (w89, w90, w88);
  c_w92     : entity work.andG  port map (w79, w80, w92);
  c_w93     : entity work.andG  port map (w78, w81, w93);
  c_w91     : entity work.orG   port map (w92, w93, w91);
  c_w87     : entity work.xorG  port map (w88, w91, w87);
  c_w96     : entity work.wire  port map (a_12, w96);
  c_w97     : entity work.wire  port map (b_12, w97);
  c_w95     : entity work.xorG  port map (w96, w97, w95);
  c_w101    : entity work.andG  port map (w89, w90, w101);
  c_w102    : entity work.andG  port map (w88, w92, w102);
  c_w100    : entity work.orG   port map (w101, w102, w100);
  c_w104    : entity work.andG  port map (w88, w78, w104);
  c_w103    : entity work.andG  port map (w104, w82, w103);
  c_w99     : entity work.orG   port map (w100, w103, w99);
  c_w106    : entity work.andG  port map (w104, w86, w106);
  c_w105    : entity work.andG  port map (w106, w61, w105);
  c_w98     : entity work.orG   port map (w99, w105, w98);
  c_w94     : entity work.xorG  port map (w95, w98, w94);
  c_w109    : entity work.wire  port map (a_13, w109);
  c_w110    : entity work.wire  port map (b_13, w110);
  c_w108    : entity work.xorG  port map (w109, w110, w108);
  c_w112    : entity work.andG  port map (w96, w97, w112);
  c_w113    : entity work.andG  port map (w95, w98, w113);
  c_w111    : entity work.orG   port map (w112, w113, w111);
  c_w107    : entity work.xorG  port map (w108, w111, w107);
  c_w116    : entity work.wire  port map (a_14, w116);
  c_w117    : entity work.wire  port map (b_14, w117);
  c_w115    : entity work.xorG  port map (w116, w117, w115);
  c_w120    : entity work.andG  port map (w109, w110, w120);
  c_w121    : entity work.andG  port map (w108, w112, w121);
  c_w119    : entity work.orG   port map (w120, w121, w119);
  c_w123    : entity work.andG  port map (w108, w95, w123);
  c_w122    : entity work.andG  port map (w123, w98, w122);
  c_w118    : entity work.orG   port map (w119, w122, w118);
  c_w114    : entity work.xorG  port map (w115, w118, w114);
  c_w126    : entity work.wire  port map (a_15, w126);
  c_w127    : entity work.wire  port map (b_15, w127);
  c_w125    : entity work.xorG  port map (w126, w127, w125);
  c_w129    : entity work.andG  port map (w116, w117, w129);
  c_w130    : entity work.andG  port map (w115, w118, w130);
  c_w128    : entity work.orG   port map (w129, w130, w128);
  c_w124    : entity work.xorG  port map (w125, w128, w124);
  c_w133    : entity work.wire  port map (a_16, w133);
  c_w134    : entity work.wire  port map (b_16, w134);
  c_w132    : entity work.xorG  port map (w133, w134, w132);
  c_w139    : entity work.andG  port map (w126, w127, w139);
  c_w140    : entity work.andG  port map (w125, w129, w140);
  c_w138    : entity work.orG   port map (w139, w140, w138);
  c_w142    : entity work.andG  port map (w125, w115, w142);
  c_w141    : entity work.andG  port map (w142, w119, w141);
  c_w137    : entity work.orG   port map (w138, w141, w137);
  c_w144    : entity work.andG  port map (w142, w123, w144);
  c_w143    : entity work.andG  port map (w144, w99, w143);
  c_w136    : entity work.orG   port map (w137, w143, w136);
  c_w146    : entity work.andG  port map (w144, w106, w146);
  c_w145    : entity work.andG  port map (w146, w61, w145);
  c_w135    : entity work.orG   port map (w136, w145, w135);
  c_w131    : entity work.xorG  port map (w132, w135, w131);
  c_w149    : entity work.wire  port map (a_17, w149);
  c_w150    : entity work.wire  port map (b_17, w150);
  c_w148    : entity work.xorG  port map (w149, w150, w148);
  c_w152    : entity work.andG  port map (w133, w134, w152);
  c_w153    : entity work.andG  port map (w132, w135, w153);
  c_w151    : entity work.orG   port map (w152, w153, w151);
  c_w147    : entity work.xorG  port map (w148, w151, w147);
  c_w156    : entity work.wire  port map (a_18, w156);
  c_w157    : entity work.wire  port map (b_18, w157);
  c_w155    : entity work.xorG  port map (w156, w157, w155);
  c_w160    : entity work.andG  port map (w149, w150, w160);
  c_w161    : entity work.andG  port map (w148, w152, w161);
  c_w159    : entity work.orG   port map (w160, w161, w159);
  c_w163    : entity work.andG  port map (w148, w132, w163);
  c_w162    : entity work.andG  port map (w163, w135, w162);
  c_w158    : entity work.orG   port map (w159, w162, w158);
  c_w154    : entity work.xorG  port map (w155, w158, w154);
  c_w166    : entity work.wire  port map (a_19, w166);
  c_w167    : entity work.wire  port map (b_19, w167);
  c_w165    : entity work.xorG  port map (w166, w167, w165);
  c_w169    : entity work.andG  port map (w156, w157, w169);
  c_w170    : entity work.andG  port map (w155, w158, w170);
  c_w168    : entity work.orG   port map (w169, w170, w168);
  c_w164    : entity work.xorG  port map (w165, w168, w164);
  c_w173    : entity work.wire  port map (a_20, w173);
  c_w174    : entity work.wire  port map (b_20, w174);
  c_w172    : entity work.xorG  port map (w173, w174, w172);
  c_w178    : entity work.andG  port map (w166, w167, w178);
  c_w179    : entity work.andG  port map (w165, w169, w179);
  c_w177    : entity work.orG   port map (w178, w179, w177);
  c_w181    : entity work.andG  port map (w165, w155, w181);
  c_w180    : entity work.andG  port map (w181, w159, w180);
  c_w176    : entity work.orG   port map (w177, w180, w176);
  c_w183    : entity work.andG  port map (w181, w163, w183);
  c_w182    : entity work.andG  port map (w183, w135, w182);
  c_w175    : entity work.orG   port map (w176, w182, w175);
  c_w171    : entity work.xorG  port map (w172, w175, w171);
  c_w186    : entity work.wire  port map (a_21, w186);
  c_w187    : entity work.wire  port map (b_21, w187);
  c_w185    : entity work.xorG  port map (w186, w187, w185);
  c_w189    : entity work.andG  port map (w173, w174, w189);
  c_w190    : entity work.andG  port map (w172, w175, w190);
  c_w188    : entity work.orG   port map (w189, w190, w188);
  c_w184    : entity work.xorG  port map (w185, w188, w184);
  c_w193    : entity work.wire  port map (a_22, w193);
  c_w194    : entity work.wire  port map (b_22, w194);
  c_w192    : entity work.xorG  port map (w193, w194, w192);
  c_w197    : entity work.andG  port map (w186, w187, w197);
  c_w198    : entity work.andG  port map (w185, w189, w198);
  c_w196    : entity work.orG   port map (w197, w198, w196);
  c_w200    : entity work.andG  port map (w185, w172, w200);
  c_w199    : entity work.andG  port map (w200, w175, w199);
  c_w195    : entity work.orG   port map (w196, w199, w195);
  c_w191    : entity work.xorG  port map (w192, w195, w191);
  c_w203    : entity work.wire  port map (a_23, w203);
  c_w204    : entity work.wire  port map (b_23, w204);
  c_w202    : entity work.xorG  port map (w203, w204, w202);
  c_w206    : entity work.andG  port map (w193, w194, w206);
  c_w207    : entity work.andG  port map (w192, w195, w207);
  c_w205    : entity work.orG   port map (w206, w207, w205);
  c_w201    : entity work.xorG  port map (w202, w205, w201);
  c_w210    : entity work.wire  port map (a_24, w210);
  c_w211    : entity work.wire  port map (b_24, w211);
  c_w209    : entity work.xorG  port map (w210, w211, w209);
  c_w216    : entity work.andG  port map (w203, w204, w216);
  c_w217    : entity work.andG  port map (w202, w206, w217);
  c_w215    : entity work.orG   port map (w216, w217, w215);
  c_w219    : entity work.andG  port map (w202, w192, w219);
  c_w218    : entity work.andG  port map (w219, w196, w218);
  c_w214    : entity work.orG   port map (w215, w218, w214);
  c_w221    : entity work.andG  port map (w219, w200, w221);
  c_w220    : entity work.andG  port map (w221, w176, w220);
  c_w213    : entity work.orG   port map (w214, w220, w213);
  c_w223    : entity work.andG  port map (w221, w183, w223);
  c_w222    : entity work.andG  port map (w223, w135, w222);
  c_w212    : entity work.orG   port map (w213, w222, w212);
  c_w208    : entity work.xorG  port map (w209, w212, w208);
  c_w226    : entity work.wire  port map (a_25, w226);
  c_w227    : entity work.wire  port map (b_25, w227);
  c_w225    : entity work.xorG  port map (w226, w227, w225);
  c_w229    : entity work.andG  port map (w210, w211, w229);
  c_w230    : entity work.andG  port map (w209, w212, w230);
  c_w228    : entity work.orG   port map (w229, w230, w228);
  c_w224    : entity work.xorG  port map (w225, w228, w224);
  c_w233    : entity work.wire  port map (a_26, w233);
  c_w234    : entity work.wire  port map (b_26, w234);
  c_w232    : entity work.xorG  port map (w233, w234, w232);
  c_w237    : entity work.andG  port map (w226, w227, w237);
  c_w238    : entity work.andG  port map (w225, w229, w238);
  c_w236    : entity work.orG   port map (w237, w238, w236);
  c_w240    : entity work.andG  port map (w225, w209, w240);
  c_w239    : entity work.andG  port map (w240, w212, w239);
  c_w235    : entity work.orG   port map (w236, w239, w235);
  c_w231    : entity work.xorG  port map (w232, w235, w231);
  c_w243    : entity work.wire  port map (a_27, w243);
  c_w244    : entity work.wire  port map (b_27, w244);
  c_w242    : entity work.xorG  port map (w243, w244, w242);
  c_w246    : entity work.andG  port map (w233, w234, w246);
  c_w247    : entity work.andG  port map (w232, w235, w247);
  c_w245    : entity work.orG   port map (w246, w247, w245);
  c_w241    : entity work.xorG  port map (w242, w245, w241);
  c_w250    : entity work.wire  port map (a_28, w250);
  c_w251    : entity work.wire  port map (b_28, w251);
  c_w249    : entity work.xorG  port map (w250, w251, w249);
  c_w255    : entity work.andG  port map (w243, w244, w255);
  c_w256    : entity work.andG  port map (w242, w246, w256);
  c_w254    : entity work.orG   port map (w255, w256, w254);
  c_w258    : entity work.andG  port map (w242, w232, w258);
  c_w257    : entity work.andG  port map (w258, w236, w257);
  c_w253    : entity work.orG   port map (w254, w257, w253);
  c_w260    : entity work.andG  port map (w258, w240, w260);
  c_w259    : entity work.andG  port map (w260, w212, w259);
  c_w252    : entity work.orG   port map (w253, w259, w252);
  c_w248    : entity work.xorG  port map (w249, w252, w248);
  c_w263    : entity work.wire  port map (a_29, w263);
  c_w264    : entity work.wire  port map (b_29, w264);
  c_w262    : entity work.xorG  port map (w263, w264, w262);
  c_w266    : entity work.andG  port map (w250, w251, w266);
  c_w267    : entity work.andG  port map (w249, w252, w267);
  c_w265    : entity work.orG   port map (w266, w267, w265);
  c_w261    : entity work.xorG  port map (w262, w265, w261);
  c_w270    : entity work.wire  port map (a_30, w270);
  c_w271    : entity work.wire  port map (b_30, w271);
  c_w269    : entity work.xorG  port map (w270, w271, w269);
  c_w274    : entity work.andG  port map (w263, w264, w274);
  c_w275    : entity work.andG  port map (w262, w266, w275);
  c_w273    : entity work.orG   port map (w274, w275, w273);
  c_w277    : entity work.andG  port map (w262, w249, w277);
  c_w276    : entity work.andG  port map (w277, w252, w276);
  c_w272    : entity work.orG   port map (w273, w276, w272);
  c_w268    : entity work.xorG  port map (w269, w272, w268);
  c_w280    : entity work.wire  port map (a_31, w280);
  c_w281    : entity work.wire  port map (b_31, w281);
  c_w279    : entity work.xorG  port map (w280, w281, w279);
  c_w283    : entity work.andG  port map (w270, w271, w283);
  c_w284    : entity work.andG  port map (w269, w272, w284);
  c_w282    : entity work.orG   port map (w283, w284, w282);
  c_w278    : entity work.xorG  port map (w279, w282, w278);
  c_w287    : entity work.wire  port map (a_32, w287);
  c_w288    : entity work.wire  port map (b_32, w288);
  c_w286    : entity work.xorG  port map (w287, w288, w286);
  c_w294    : entity work.andG  port map (w280, w281, w294);
  c_w295    : entity work.andG  port map (w279, w283, w295);
  c_w293    : entity work.orG   port map (w294, w295, w293);
  c_w297    : entity work.andG  port map (w279, w269, w297);
  c_w296    : entity work.andG  port map (w297, w273, w296);
  c_w292    : entity work.orG   port map (w293, w296, w292);
  c_w299    : entity work.andG  port map (w297, w277, w299);
  c_w298    : entity work.andG  port map (w299, w253, w298);
  c_w291    : entity work.orG   port map (w292, w298, w291);
  c_w301    : entity work.andG  port map (w299, w260, w301);
  c_w300    : entity work.andG  port map (w301, w213, w300);
  c_w290    : entity work.orG   port map (w291, w300, w290);
  c_w303    : entity work.andG  port map (w301, w223, w303);
  c_w302    : entity work.andG  port map (w303, w135, w302);
  c_w289    : entity work.orG   port map (w290, w302, w289);
  c_w285    : entity work.xorG  port map (w286, w289, w285);
  c_w306    : entity work.wire  port map (a_33, w306);
  c_w307    : entity work.wire  port map (b_33, w307);
  c_w305    : entity work.xorG  port map (w306, w307, w305);
  c_w309    : entity work.andG  port map (w287, w288, w309);
  c_w310    : entity work.andG  port map (w286, w289, w310);
  c_w308    : entity work.orG   port map (w309, w310, w308);
  c_w304    : entity work.xorG  port map (w305, w308, w304);
  c_w313    : entity work.wire  port map (a_34, w313);
  c_w314    : entity work.wire  port map (b_34, w314);
  c_w312    : entity work.xorG  port map (w313, w314, w312);
  c_w317    : entity work.andG  port map (w306, w307, w317);
  c_w318    : entity work.andG  port map (w305, w309, w318);
  c_w316    : entity work.orG   port map (w317, w318, w316);
  c_w320    : entity work.andG  port map (w305, w286, w320);
  c_w319    : entity work.andG  port map (w320, w289, w319);
  c_w315    : entity work.orG   port map (w316, w319, w315);
  c_w311    : entity work.xorG  port map (w312, w315, w311);
  c_w323    : entity work.wire  port map (a_35, w323);
  c_w324    : entity work.wire  port map (b_35, w324);
  c_w322    : entity work.xorG  port map (w323, w324, w322);
  c_w326    : entity work.andG  port map (w313, w314, w326);
  c_w327    : entity work.andG  port map (w312, w315, w327);
  c_w325    : entity work.orG   port map (w326, w327, w325);
  c_w321    : entity work.xorG  port map (w322, w325, w321);
  c_w330    : entity work.wire  port map (a_36, w330);
  c_w331    : entity work.wire  port map (b_36, w331);
  c_w329    : entity work.xorG  port map (w330, w331, w329);
  c_w335    : entity work.andG  port map (w323, w324, w335);
  c_w336    : entity work.andG  port map (w322, w326, w336);
  c_w334    : entity work.orG   port map (w335, w336, w334);
  c_w338    : entity work.andG  port map (w322, w312, w338);
  c_w337    : entity work.andG  port map (w338, w316, w337);
  c_w333    : entity work.orG   port map (w334, w337, w333);
  c_w340    : entity work.andG  port map (w338, w320, w340);
  c_w339    : entity work.andG  port map (w340, w289, w339);
  c_w332    : entity work.orG   port map (w333, w339, w332);
  c_w328    : entity work.xorG  port map (w329, w332, w328);
  c_w343    : entity work.wire  port map (a_37, w343);
  c_w344    : entity work.wire  port map (b_37, w344);
  c_w342    : entity work.xorG  port map (w343, w344, w342);
  c_w346    : entity work.andG  port map (w330, w331, w346);
  c_w347    : entity work.andG  port map (w329, w332, w347);
  c_w345    : entity work.orG   port map (w346, w347, w345);
  c_w341    : entity work.xorG  port map (w342, w345, w341);
  c_w350    : entity work.wire  port map (a_38, w350);
  c_w351    : entity work.wire  port map (b_38, w351);
  c_w349    : entity work.xorG  port map (w350, w351, w349);
  c_w354    : entity work.andG  port map (w343, w344, w354);
  c_w355    : entity work.andG  port map (w342, w346, w355);
  c_w353    : entity work.orG   port map (w354, w355, w353);
  c_w357    : entity work.andG  port map (w342, w329, w357);
  c_w356    : entity work.andG  port map (w357, w332, w356);
  c_w352    : entity work.orG   port map (w353, w356, w352);
  c_w348    : entity work.xorG  port map (w349, w352, w348);
  c_w360    : entity work.wire  port map (a_39, w360);
  c_w361    : entity work.wire  port map (b_39, w361);
  c_w359    : entity work.xorG  port map (w360, w361, w359);
  c_w363    : entity work.andG  port map (w350, w351, w363);
  c_w364    : entity work.andG  port map (w349, w352, w364);
  c_w362    : entity work.orG   port map (w363, w364, w362);
  c_w358    : entity work.xorG  port map (w359, w362, w358);
  c_w367    : entity work.wire  port map (a_40, w367);
  c_w368    : entity work.wire  port map (b_40, w368);
  c_w366    : entity work.xorG  port map (w367, w368, w366);
  c_w373    : entity work.andG  port map (w360, w361, w373);
  c_w374    : entity work.andG  port map (w359, w363, w374);
  c_w372    : entity work.orG   port map (w373, w374, w372);
  c_w376    : entity work.andG  port map (w359, w349, w376);
  c_w375    : entity work.andG  port map (w376, w353, w375);
  c_w371    : entity work.orG   port map (w372, w375, w371);
  c_w378    : entity work.andG  port map (w376, w357, w378);
  c_w377    : entity work.andG  port map (w378, w333, w377);
  c_w370    : entity work.orG   port map (w371, w377, w370);
  c_w380    : entity work.andG  port map (w378, w340, w380);
  c_w379    : entity work.andG  port map (w380, w289, w379);
  c_w369    : entity work.orG   port map (w370, w379, w369);
  c_w365    : entity work.xorG  port map (w366, w369, w365);
  c_w383    : entity work.wire  port map (a_41, w383);
  c_w384    : entity work.wire  port map (b_41, w384);
  c_w382    : entity work.xorG  port map (w383, w384, w382);
  c_w386    : entity work.andG  port map (w367, w368, w386);
  c_w387    : entity work.andG  port map (w366, w369, w387);
  c_w385    : entity work.orG   port map (w386, w387, w385);
  c_w381    : entity work.xorG  port map (w382, w385, w381);
  c_w390    : entity work.wire  port map (a_42, w390);
  c_w391    : entity work.wire  port map (b_42, w391);
  c_w389    : entity work.xorG  port map (w390, w391, w389);
  c_w394    : entity work.andG  port map (w383, w384, w394);
  c_w395    : entity work.andG  port map (w382, w386, w395);
  c_w393    : entity work.orG   port map (w394, w395, w393);
  c_w397    : entity work.andG  port map (w382, w366, w397);
  c_w396    : entity work.andG  port map (w397, w369, w396);
  c_w392    : entity work.orG   port map (w393, w396, w392);
  c_w388    : entity work.xorG  port map (w389, w392, w388);
  c_w400    : entity work.wire  port map (a_43, w400);
  c_w401    : entity work.wire  port map (b_43, w401);
  c_w399    : entity work.xorG  port map (w400, w401, w399);
  c_w403    : entity work.andG  port map (w390, w391, w403);
  c_w404    : entity work.andG  port map (w389, w392, w404);
  c_w402    : entity work.orG   port map (w403, w404, w402);
  c_w398    : entity work.xorG  port map (w399, w402, w398);
  c_w407    : entity work.wire  port map (a_44, w407);
  c_w408    : entity work.wire  port map (b_44, w408);
  c_w406    : entity work.xorG  port map (w407, w408, w406);
  c_w412    : entity work.andG  port map (w400, w401, w412);
  c_w413    : entity work.andG  port map (w399, w403, w413);
  c_w411    : entity work.orG   port map (w412, w413, w411);
  c_w415    : entity work.andG  port map (w399, w389, w415);
  c_w414    : entity work.andG  port map (w415, w393, w414);
  c_w410    : entity work.orG   port map (w411, w414, w410);
  c_w417    : entity work.andG  port map (w415, w397, w417);
  c_w416    : entity work.andG  port map (w417, w369, w416);
  c_w409    : entity work.orG   port map (w410, w416, w409);
  c_w405    : entity work.xorG  port map (w406, w409, w405);
  c_w420    : entity work.wire  port map (a_45, w420);
  c_w421    : entity work.wire  port map (b_45, w421);
  c_w419    : entity work.xorG  port map (w420, w421, w419);
  c_w423    : entity work.andG  port map (w407, w408, w423);
  c_w424    : entity work.andG  port map (w406, w409, w424);
  c_w422    : entity work.orG   port map (w423, w424, w422);
  c_w418    : entity work.xorG  port map (w419, w422, w418);
  c_w427    : entity work.wire  port map (a_46, w427);
  c_w428    : entity work.wire  port map (b_46, w428);
  c_w426    : entity work.xorG  port map (w427, w428, w426);
  c_w431    : entity work.andG  port map (w420, w421, w431);
  c_w432    : entity work.andG  port map (w419, w423, w432);
  c_w430    : entity work.orG   port map (w431, w432, w430);
  c_w434    : entity work.andG  port map (w419, w406, w434);
  c_w433    : entity work.andG  port map (w434, w409, w433);
  c_w429    : entity work.orG   port map (w430, w433, w429);
  c_w425    : entity work.xorG  port map (w426, w429, w425);
  c_w437    : entity work.wire  port map (a_47, w437);
  c_w438    : entity work.wire  port map (b_47, w438);
  c_w436    : entity work.xorG  port map (w437, w438, w436);
  c_w440    : entity work.andG  port map (w427, w428, w440);
  c_w441    : entity work.andG  port map (w426, w429, w441);
  c_w439    : entity work.orG   port map (w440, w441, w439);
  c_w435    : entity work.xorG  port map (w436, w439, w435);
  c_w444    : entity work.wire  port map (a_48, w444);
  c_w445    : entity work.wire  port map (b_48, w445);
  c_w443    : entity work.xorG  port map (w444, w445, w443);
  c_w451    : entity work.andG  port map (w437, w438, w451);
  c_w452    : entity work.andG  port map (w436, w440, w452);
  c_w450    : entity work.orG   port map (w451, w452, w450);
  c_w454    : entity work.andG  port map (w436, w426, w454);
  c_w453    : entity work.andG  port map (w454, w430, w453);
  c_w449    : entity work.orG   port map (w450, w453, w449);
  c_w456    : entity work.andG  port map (w454, w434, w456);
  c_w455    : entity work.andG  port map (w456, w410, w455);
  c_w448    : entity work.orG   port map (w449, w455, w448);
  c_w458    : entity work.andG  port map (w456, w417, w458);
  c_w457    : entity work.andG  port map (w458, w370, w457);
  c_w447    : entity work.orG   port map (w448, w457, w447);
  c_w460    : entity work.andG  port map (w458, w380, w460);
  c_w459    : entity work.andG  port map (w460, w289, w459);
  c_w446    : entity work.orG   port map (w447, w459, w446);
  c_w442    : entity work.xorG  port map (w443, w446, w442);
  c_w463    : entity work.wire  port map (a_49, w463);
  c_w464    : entity work.wire  port map (b_49, w464);
  c_w462    : entity work.xorG  port map (w463, w464, w462);
  c_w466    : entity work.andG  port map (w444, w445, w466);
  c_w467    : entity work.andG  port map (w443, w446, w467);
  c_w465    : entity work.orG   port map (w466, w467, w465);
  c_w461    : entity work.xorG  port map (w462, w465, w461);
  c_w470    : entity work.wire  port map (a_50, w470);
  c_w471    : entity work.wire  port map (b_50, w471);
  c_w469    : entity work.xorG  port map (w470, w471, w469);
  c_w474    : entity work.andG  port map (w463, w464, w474);
  c_w475    : entity work.andG  port map (w462, w466, w475);
  c_w473    : entity work.orG   port map (w474, w475, w473);
  c_w477    : entity work.andG  port map (w462, w443, w477);
  c_w476    : entity work.andG  port map (w477, w446, w476);
  c_w472    : entity work.orG   port map (w473, w476, w472);
  c_w468    : entity work.xorG  port map (w469, w472, w468);
  c_w480    : entity work.wire  port map (a_51, w480);
  c_w481    : entity work.wire  port map (b_51, w481);
  c_w479    : entity work.xorG  port map (w480, w481, w479);
  c_w483    : entity work.andG  port map (w470, w471, w483);
  c_w484    : entity work.andG  port map (w469, w472, w484);
  c_w482    : entity work.orG   port map (w483, w484, w482);
  c_w478    : entity work.xorG  port map (w479, w482, w478);
  c_w487    : entity work.wire  port map (a_52, w487);
  c_w488    : entity work.wire  port map (b_52, w488);
  c_w486    : entity work.xorG  port map (w487, w488, w486);
  c_w492    : entity work.andG  port map (w480, w481, w492);
  c_w493    : entity work.andG  port map (w479, w483, w493);
  c_w491    : entity work.orG   port map (w492, w493, w491);
  c_w495    : entity work.andG  port map (w479, w469, w495);
  c_w494    : entity work.andG  port map (w495, w473, w494);
  c_w490    : entity work.orG   port map (w491, w494, w490);
  c_w497    : entity work.andG  port map (w495, w477, w497);
  c_w496    : entity work.andG  port map (w497, w446, w496);
  c_w489    : entity work.orG   port map (w490, w496, w489);
  c_w485    : entity work.xorG  port map (w486, w489, w485);
  c_w500    : entity work.wire  port map (a_53, w500);
  c_w501    : entity work.wire  port map (b_53, w501);
  c_w499    : entity work.xorG  port map (w500, w501, w499);
  c_w503    : entity work.andG  port map (w487, w488, w503);
  c_w504    : entity work.andG  port map (w486, w489, w504);
  c_w502    : entity work.orG   port map (w503, w504, w502);
  c_w498    : entity work.xorG  port map (w499, w502, w498);
  c_w507    : entity work.wire  port map (a_54, w507);
  c_w508    : entity work.wire  port map (b_54, w508);
  c_w506    : entity work.xorG  port map (w507, w508, w506);
  c_w511    : entity work.andG  port map (w500, w501, w511);
  c_w512    : entity work.andG  port map (w499, w503, w512);
  c_w510    : entity work.orG   port map (w511, w512, w510);
  c_w514    : entity work.andG  port map (w499, w486, w514);
  c_w513    : entity work.andG  port map (w514, w489, w513);
  c_w509    : entity work.orG   port map (w510, w513, w509);
  c_w505    : entity work.xorG  port map (w506, w509, w505);
  c_w517    : entity work.wire  port map (a_55, w517);
  c_w518    : entity work.wire  port map (b_55, w518);
  c_w516    : entity work.xorG  port map (w517, w518, w516);
  c_w520    : entity work.andG  port map (w507, w508, w520);
  c_w521    : entity work.andG  port map (w506, w509, w521);
  c_w519    : entity work.orG   port map (w520, w521, w519);
  c_w515    : entity work.xorG  port map (w516, w519, w515);
  c_w524    : entity work.wire  port map (a_56, w524);
  c_w525    : entity work.wire  port map (b_56, w525);
  c_w523    : entity work.xorG  port map (w524, w525, w523);
  c_w530    : entity work.andG  port map (w517, w518, w530);
  c_w531    : entity work.andG  port map (w516, w520, w531);
  c_w529    : entity work.orG   port map (w530, w531, w529);
  c_w533    : entity work.andG  port map (w516, w506, w533);
  c_w532    : entity work.andG  port map (w533, w510, w532);
  c_w528    : entity work.orG   port map (w529, w532, w528);
  c_w535    : entity work.andG  port map (w533, w514, w535);
  c_w534    : entity work.andG  port map (w535, w490, w534);
  c_w527    : entity work.orG   port map (w528, w534, w527);
  c_w537    : entity work.andG  port map (w535, w497, w537);
  c_w536    : entity work.andG  port map (w537, w446, w536);
  c_w526    : entity work.orG   port map (w527, w536, w526);
  c_w522    : entity work.xorG  port map (w523, w526, w522);
  c_w540    : entity work.wire  port map (a_57, w540);
  c_w541    : entity work.wire  port map (b_57, w541);
  c_w539    : entity work.xorG  port map (w540, w541, w539);
  c_w543    : entity work.andG  port map (w524, w525, w543);
  c_w544    : entity work.andG  port map (w523, w526, w544);
  c_w542    : entity work.orG   port map (w543, w544, w542);
  c_w538    : entity work.xorG  port map (w539, w542, w538);
  c_w547    : entity work.wire  port map (a_58, w547);
  c_w548    : entity work.wire  port map (b_58, w548);
  c_w546    : entity work.xorG  port map (w547, w548, w546);
  c_w551    : entity work.andG  port map (w540, w541, w551);
  c_w552    : entity work.andG  port map (w539, w543, w552);
  c_w550    : entity work.orG   port map (w551, w552, w550);
  c_w554    : entity work.andG  port map (w539, w523, w554);
  c_w553    : entity work.andG  port map (w554, w526, w553);
  c_w549    : entity work.orG   port map (w550, w553, w549);
  c_w545    : entity work.xorG  port map (w546, w549, w545);
  c_w557    : entity work.wire  port map (a_59, w557);
  c_w558    : entity work.wire  port map (b_59, w558);
  c_w556    : entity work.xorG  port map (w557, w558, w556);
  c_w560    : entity work.andG  port map (w547, w548, w560);
  c_w561    : entity work.andG  port map (w546, w549, w561);
  c_w559    : entity work.orG   port map (w560, w561, w559);
  c_w555    : entity work.xorG  port map (w556, w559, w555);
  c_w564    : entity work.wire  port map (a_60, w564);
  c_w565    : entity work.wire  port map (b_60, w565);
  c_w563    : entity work.xorG  port map (w564, w565, w563);
  c_w569    : entity work.andG  port map (w557, w558, w569);
  c_w570    : entity work.andG  port map (w556, w560, w570);
  c_w568    : entity work.orG   port map (w569, w570, w568);
  c_w572    : entity work.andG  port map (w556, w546, w572);
  c_w571    : entity work.andG  port map (w572, w550, w571);
  c_w567    : entity work.orG   port map (w568, w571, w567);
  c_w574    : entity work.andG  port map (w572, w554, w574);
  c_w573    : entity work.andG  port map (w574, w526, w573);
  c_w566    : entity work.orG   port map (w567, w573, w566);
  c_w562    : entity work.xorG  port map (w563, w566, w562);
  c_w577    : entity work.wire  port map (a_61, w577);
  c_w578    : entity work.wire  port map (b_61, w578);
  c_w576    : entity work.xorG  port map (w577, w578, w576);
  c_w580    : entity work.andG  port map (w564, w565, w580);
  c_w581    : entity work.andG  port map (w563, w566, w581);
  c_w579    : entity work.orG   port map (w580, w581, w579);
  c_w575    : entity work.xorG  port map (w576, w579, w575);
  c_w584    : entity work.wire  port map (a_62, w584);
  c_w585    : entity work.wire  port map (b_62, w585);
  c_w583    : entity work.xorG  port map (w584, w585, w583);
  c_w588    : entity work.andG  port map (w577, w578, w588);
  c_w589    : entity work.andG  port map (w576, w580, w589);
  c_w587    : entity work.orG   port map (w588, w589, w587);
  c_w591    : entity work.andG  port map (w576, w563, w591);
  c_w590    : entity work.andG  port map (w591, w566, w590);
  c_w586    : entity work.orG   port map (w587, w590, w586);
  c_w582    : entity work.xorG  port map (w583, w586, w582);
  c_w594    : entity work.wire  port map (a_63, w594);
  c_w595    : entity work.wire  port map (b_63, w595);
  c_w593    : entity work.xorG  port map (w594, w595, w593);
  c_w597    : entity work.andG  port map (w584, w585, w597);
  c_w598    : entity work.andG  port map (w583, w586, w598);
  c_w596    : entity work.orG   port map (w597, w598, w596);
  c_w592    : entity work.xorG  port map (w593, w596, w592);
  c_w605    : entity work.andG  port map (w594, w595, w605);
  c_w606    : entity work.andG  port map (w593, w597, w606);
  c_w604    : entity work.orG   port map (w605, w606, w604);
  c_w608    : entity work.andG  port map (w593, w583, w608);
  c_w607    : entity work.andG  port map (w608, w587, w607);
  c_w603    : entity work.orG   port map (w604, w607, w603);
  c_w610    : entity work.andG  port map (w608, w591, w610);
  c_w609    : entity work.andG  port map (w610, w567, w609);
  c_w602    : entity work.orG   port map (w603, w609, w602);
  c_w612    : entity work.andG  port map (w610, w574, w612);
  c_w611    : entity work.andG  port map (w612, w527, w611);
  c_w601    : entity work.orG   port map (w602, w611, w601);
  c_w614    : entity work.andG  port map (w612, w537, w614);
  c_w613    : entity work.andG  port map (w614, w447, w613);
  c_w600    : entity work.orG   port map (w601, w613, w600);
  c_w616    : entity work.andG  port map (w614, w460, w616);
  c_w615    : entity work.andG  port map (w616, w289, w615);
  c_w599    : entity work.orG   port map (w600, w615, w599);

  
  c_sum_0   : entity work.wire  port map (w1, sum_0);
  c_sum_1   : entity work.wire  port map (w4, sum_1);
  c_sum_2   : entity work.wire  port map (w9, sum_2);
  c_sum_3   : entity work.wire  port map (w16, sum_3);
  c_sum_4   : entity work.wire  port map (w23, sum_4);
  c_sum_5   : entity work.wire  port map (w33, sum_5);
  c_sum_6   : entity work.wire  port map (w40, sum_6);
  c_sum_7   : entity work.wire  port map (w50, sum_7);
  c_sum_8   : entity work.wire  port map (w57, sum_8);
  c_sum_9   : entity work.wire  port map (w70, sum_9);
  c_sum_10  : entity work.wire  port map (w77, sum_10);
  c_sum_11  : entity work.wire  port map (w87, sum_11);
  c_sum_12  : entity work.wire  port map (w94, sum_12);
  c_sum_13  : entity work.wire  port map (w107, sum_13);
  c_sum_14  : entity work.wire  port map (w114, sum_14);
  c_sum_15  : entity work.wire  port map (w124, sum_15);
  c_sum_16  : entity work.wire  port map (w131, sum_16);
  c_sum_17  : entity work.wire  port map (w147, sum_17);
  c_sum_18  : entity work.wire  port map (w154, sum_18);
  c_sum_19  : entity work.wire  port map (w164, sum_19);
  c_sum_20  : entity work.wire  port map (w171, sum_20);
  c_sum_21  : entity work.wire  port map (w184, sum_21);
  c_sum_22  : entity work.wire  port map (w191, sum_22);
  c_sum_23  : entity work.wire  port map (w201, sum_23);
  c_sum_24  : entity work.wire  port map (w208, sum_24);
  c_sum_25  : entity work.wire  port map (w224, sum_25);
  c_sum_26  : entity work.wire  port map (w231, sum_26);
  c_sum_27  : entity work.wire  port map (w241, sum_27);
  c_sum_28  : entity work.wire  port map (w248, sum_28);
  c_sum_29  : entity work.wire  port map (w261, sum_29);
  c_sum_30  : entity work.wire  port map (w268, sum_30);
  c_sum_31  : entity work.wire  port map (w278, sum_31);
  c_sum_32  : entity work.wire  port map (w285, sum_32);
  c_sum_33  : entity work.wire  port map (w304, sum_33);
  c_sum_34  : entity work.wire  port map (w311, sum_34);
  c_sum_35  : entity work.wire  port map (w321, sum_35);
  c_sum_36  : entity work.wire  port map (w328, sum_36);
  c_sum_37  : entity work.wire  port map (w341, sum_37);
  c_sum_38  : entity work.wire  port map (w348, sum_38);
  c_sum_39  : entity work.wire  port map (w358, sum_39);
  c_sum_40  : entity work.wire  port map (w365, sum_40);
  c_sum_41  : entity work.wire  port map (w381, sum_41);
  c_sum_42  : entity work.wire  port map (w388, sum_42);
  c_sum_43  : entity work.wire  port map (w398, sum_43);
  c_sum_44  : entity work.wire  port map (w405, sum_44);
  c_sum_45  : entity work.wire  port map (w418, sum_45);
  c_sum_46  : entity work.wire  port map (w425, sum_46);
  c_sum_47  : entity work.wire  port map (w435, sum_47);
  c_sum_48  : entity work.wire  port map (w442, sum_48);
  c_sum_49  : entity work.wire  port map (w461, sum_49);
  c_sum_50  : entity work.wire  port map (w468, sum_50);
  c_sum_51  : entity work.wire  port map (w478, sum_51);
  c_sum_52  : entity work.wire  port map (w485, sum_52);
  c_sum_53  : entity work.wire  port map (w498, sum_53);
  c_sum_54  : entity work.wire  port map (w505, sum_54);
  c_sum_55  : entity work.wire  port map (w515, sum_55);
  c_sum_56  : entity work.wire  port map (w522, sum_56);
  c_sum_57  : entity work.wire  port map (w538, sum_57);
  c_sum_58  : entity work.wire  port map (w545, sum_58);
  c_sum_59  : entity work.wire  port map (w555, sum_59);
  c_sum_60  : entity work.wire  port map (w562, sum_60);
  c_sum_61  : entity work.wire  port map (w575, sum_61);
  c_sum_62  : entity work.wire  port map (w582, sum_62);
  c_sum_63  : entity work.wire  port map (w592, sum_63);
  c_cout    : entity work.wire  port map (w599, cout);
end structural;
